library ieee;
use ieee.std_logic_1164.all;

package common_p is
	type logic_matrix_t is array(natural range <>, natural range<>) of std_logic;
end common_p;

package body common_p is
end common_p;